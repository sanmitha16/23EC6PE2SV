interface atm_if;
    logic clk;
    logic reset;
    logic card_inserted;
    logic pin_correct;
    logic balance_ok;
    logic dispense_cash;
endinterface
interface atm_if;
    logic clk;
    logic reset;
    logic card_inserted;
    logic pin_correct;
    logic balance_ok;
    logic dispense_cash;
endinterface